`timescale 1ns / 1ps

module test_spi
(
    inout wire sclk,
    inout wire mosi,
    inout wire miso,
    inout wire ncs,
    inout wire [1:0] spi_mode,
    inout wire [5:0] spi_word_width
);

endmodule // test_spi
