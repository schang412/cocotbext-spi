`timescale 1ns / 1ps

module test_tmc4671
(
    inout wire sclk,
    inout wire mosi,
    inout wire miso,
    inout wire ncs
);

endmodule // test_tmc4671
