`timescale 1ns / 1ps

module test_drv8304
(
    inout wire sclk,
    inout wire mosi,
    inout wire miso,
    inout wire ncs
);

endmodule // test_drv8304
