`timescale 1ns / 1ps

module test_ads8028
(
    inout wire sclk,
    inout wire mosi,
    inout wire miso,
    inout wire ncs
);

endmodule // test_ads8028